package ram_pkg;
	// import uvm_pkg
   	import uvm_pkg::*;

	// include the uvm_macros.svh
    `include "uvm_macros.svh"

  
	// include the tb_defs.sv
    `include "tb_defs.sv"

 	//include write_xtn.sv  
    `include "write_xtn.sv"  

endpackage
